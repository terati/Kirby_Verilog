//NVM