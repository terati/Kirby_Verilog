

  
//-------------------------------------------------------------------------
//      VGA controller                                                   --
//      Kyle Kloepper                                                    --
//      4-05-2005                                                        --
//                                                                       --
//      Modified by Stephen Kempf 04-08-2005                             --
//                                10-05-2006                             --
//                                03-12-2007                             --
//      Translated by Joe Meng    07-07-2013                             --
//      Modified by Po-Han Huang  12-08-2017                             --
//      Spring 2018 Distribution                                         --
//                                                                       --
//      Used standard 640x480 vga found at epanorama                     --
//                                                                       --
//      reference: http://www.xilinx.com/bvdocs/userguides/ug130.pdf     --
//                 http://www.epanorama.net/documents/pc/vga_timing.html --
//                                                                       -- 
//      note: The standard is changed slightly because of 25 mhz instead --
//            of 25.175 mhz pixel clock. Refresh rate drops slightly.    --
//                                                                       --
//      For use with ECE 385 Lab 8 and Final Project                     --
//      ECE Department @ UIUC                                            --
//-------------------------------------------------------------------------


module  VGA_controller (input              Clk,         // 50 MHz clock
                                           Reset,       // Active-high reset signal
														 FAST_CLK,	  // 100 MHz clock
														 BOSSTIME,
                        output logic       VGA_HS,      // Horizontal sync pulse.  Active low
                                           VGA_VS,      // Vertical sync pulse.  Active low
                        input             VGA_CLK,     // 25 MHz VGA clock input
                        output logic       VGA_BLANK_N, // Blanking interval indicator.  Active low.
                                           VGA_SYNC_N,  // Composite Sync signal.  Active low.  We don't use it in this lab,
                                                        // but the video DAC on the DE2 board requires an input for it.
                        output logic [9:0] DrawX,       // horizontal coordinate
                                           DrawY,       // vertical coordinate
												
								output logic [7:0] VGA_R, VGA_G, VGA_B, 
								input logic		 is_kirby_temp, is_block_temp, is_waddle0_temp, is_attack_temp, is_background_temp, is_atk_temp, boss, is_flame,
								output logic 		 is_kirby, is_block, is_attack, is_background,
								input logic [7:0]  Red, Green, Blue, kred, kgreen, kblue, wred, wgreen, wblue, kirbydata, atkdata, ared, agreen, ablue, bred, bgreen, bblue, Batkdata, waddledata
								
                        );     
    
    // 800 pixels per line (including front/back porch)
    // 525 lines per frame (including front/back porch)
    parameter [9:0] H_TOTAL = 10'd800;
    parameter [9:0] V_TOTAL = 10'd525;
    
    logic VGA_HS_in, VGA_VS_in, VGA_BLANK_N_in, background_compare, attack_compare, block_compare, kirby_compare;
    logic [9:0] h_counter, v_counter;
    logic [9:0] h_counter_in, v_counter_in;
	 logic [7:0] red_attack_temp, blue_attack_temp, green_attack_temp, red_kirby_temp, blue_kirby_temp, green_kirby_temp,
	 red_block_temp, green_block_temp, blue_block_temp, red_background_temp, green_background_temp, blue_background_temp;
	 logic [7:0] VGA_R_temp, VGA_G_temp, VGA_B_temp;
   

	
    assign VGA_SYNC_N = 1'b0;
    assign DrawX = h_counter;
    assign DrawY = v_counter;

	 logic [1:0] State = 2'd0;
    localparam ATTACK         = 2'd0;
    localparam KIRBY          = 2'd1;
    localparam ENEMY_BLOCK    = 2'd2;
    localparam BACKGROUND     = 2'd3;
    
    // VGA control signals. 
    // VGA_CLK is generated by PLL, so you will have to manually generate it in simulation.
    always_ff @ (posedge VGA_CLK)
    begin
				if (Reset)
				  begin
						VGA_HS <= 1'b0;
						VGA_VS <= 1'b0;
						VGA_BLANK_N <= 1'b0;
						h_counter <= 10'd0;
						v_counter <= 10'd0;
				  end
				  else
				  begin
						VGA_HS <= VGA_HS_in;
						VGA_VS <= VGA_VS_in;
						VGA_BLANK_N <= VGA_BLANK_N_in;
						h_counter <= h_counter_in;
						v_counter <= v_counter_in;
				  end
				  
				  case(State)
						2'd0: begin
							is_kirby <= 1'b0; 
							is_block <= 1'b1;
							is_attack <= 1'b0;
							if(BOSSTIME) begin
								State <= State + 1;
							end
						end
						
						2'd1: begin
							is_kirby <= 1'b1; 
							is_block <= 1'b0;
							is_attack <= 1'b0;
						end
					endcase
    end

    
    always_comb
    begin
        // horizontal and vertical counter
        h_counter_in = h_counter + 10'd1;
        v_counter_in = v_counter;
        if(h_counter + 10'd1 == H_TOTAL)
        begin
            h_counter_in = 10'd0;
            if(v_counter + 10'd1 == V_TOTAL)
                v_counter_in = 10'd0;
            else
                v_counter_in = v_counter + 10'd1;
        end
        // Horizontal sync pulse is 96 pixels long at pixels 656-752
        // (Signal is registered to ensure clean output waveform)
        VGA_HS_in = 1'b1;
        if(h_counter_in >= 10'd656 && h_counter_in < 10'd752)
            VGA_HS_in = 1'b0;
        // Vertical sync pulse is 2 lines (800 pixels each) long at line 490-491
        //(Signal is registered to ensure clean output waveform)
        VGA_VS_in = 1'b1;
        if(v_counter_in >= 10'd490 && v_counter_in < 10'd492)
            VGA_VS_in = 1'b0;
        // Display pixels (inhibit blanking) between horizontal 0-639 and vertical 0-479 (640x480)
        VGA_BLANK_N_in = 1'b0;
        if(h_counter_in < 10'd640 && v_counter_in < 10'd480)
            VGA_BLANK_N_in = 1'b1;
				
				
		  VGA_R = Red;
		  VGA_G = Green;
		  VGA_B = Blue;
		  
		 
		  if((waddledata != 8'b111010)  && (is_waddle0_temp)) begin  //waddle
			  VGA_R = wred;
			  VGA_G = wgreen;
			  VGA_B = wblue;
		  end  
		  
		  if((Batkdata != 8'b111010) && (is_flame)) begin
			  VGA_R = bred;
			  VGA_G = bgreen;
			  VGA_B = bblue;
		  end 
		  
		  if((waddledata != 8'b111010) && (boss)) begin
			  VGA_R = wred;
			  VGA_G = wgreen;
			  VGA_B = wblue;
		  end 
		  
		  if((atkdata != 8'b111010) && (is_atk_temp)) begin			//atk
			  VGA_R = ared;
			  VGA_G = agreen;
			  VGA_B = ablue;
		  end 
		  
		  if((kirbydata != 8'b111010) && (is_kirby_temp)) begin	//kirby
			  VGA_R = kred;
			  VGA_G = kgreen;
			  VGA_B = kblue;
		  end 
		    
		  
		  
    end
    
endmodule

