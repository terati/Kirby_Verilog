//nvm bruh